import uarch_pkg::*;