module alu_rs
import riscv_isa_pkg::*; 
import uarch_pkg::*;
 #(
    RS_SIZE = 5
 )(
   //wip
    input logic clk, rst, flush, cache_stall,
    // Ports from Displatch
    input instruction_t rs_entry[PIPE_WIDTH - 1 : 0],

    input logic [PIPE_WIDTH - 1 : 0] rs_we,
    //Ports to Dispatch
    output logic [PIPE_WIDTH - 1 : 0] rs_rdy, //2,1,0 = 2+, 1, 0
    //Ports to Execute
    output  instruction_t execute_pkt [1:0],
    //Ports from Execute
    input logic [1:0] alu_rdy,
    //CDB PORT 
    input writeback_packet_t cdb_ports [PIPE_WIDTH - 1 : 0] 
);
//how many alu we have
function int oh_2_i (logic [PIPE_WIDTH-1:0] v);
        int o;
        o = -1;
        for (int i = 0; i < PIPE_WIDTH; i++) if (v[i]) o = i;
        return o;
    endfunction


logic [RS_SIZE - 1 : 0] indv_rs_we;
logic [RS_SIZE - 1 : 0] indv_rs_write_rdy ;
logic [RS_SIZE - 1 : 0] [PIPE_WIDTH - 1 : 0]  rs_sel;
logic [RS_SIZE - 1 : 0] indv_rs_read_rdy ;
logic [RS_SIZE - 1 : 0] indv_alu_rdy ;
instruction_t indv_execute_pkt [RS_SIZE - 1 : 0];
instruction_t muxed_rs_entry [RS_SIZE - 1 : 0];

genvar i;
generate
    for (i = 0; i < RS_SIZE; i++) begin
        rs rs(
        .clk(clk), 
        .rst(rst), 
        .flush(flush), 
        .cache_stall(cache_stall),
        // Ports from Displatch
        .rs_entry(muxed_rs_entry[i]),
        .rs_we(indv_rs_we[i]),
        //Ports to Dispatch
        .rs_write_rdy(indv_rs_write_rdy[i]),
        .rs_read_rdy(indv_rs_read_rdy[i]),
        //Ports to Execute
        .execute_pkt(indv_execute_pkt[i]),
        //Ports from Execute
        .alu_re(indv_alu_rdy[i]),
        //CDB PORT 
        .cdb_ports(cdb_ports));
    end

endgenerate

logic [$clog2(PIPE_WIDTH) + 1 : 0] s;
logic [$clog2(RS_SIZE) + 1 : 0] total_open_entries, total_ready_entries;
function int ret_exe_candidate(int best_no);
    instruction_t candidate [RS_SIZE];
    int o [RS_SIZE];
    foreach(candidate[i]) candidate[i] = '0;

    for(int i = 0; i < best_no; i++) begin
        foreach(indv_execute_pkt[j]) begin
            if(indv_rs_read_rdy[j]) begin
                if(candidate[i] == '0)begin
                     candidate[i] = indv_execute_pkt[j];
                     o[i] = j;
                end
                else if (indv_execute_pkt[j].pc < candidate[i].pc)begin
                    if(i == 0) begin
                        candidate[i] = indv_execute_pkt[j];
                        o[i] = j;
                    end
                    else if (o[i] != o[i - 1]) begin
                        candidate[i] = indv_execute_pkt[j];
                        o[i] = j;
                    end
                end
            end
        end
    end
    return o[best_no - 1];
endfunction

int c1, c2;
always_comb begin
    s = 0;
    foreach (indv_alu_rdy[i]) indv_alu_rdy[i] = 1'b0;
    total_open_entries = '0;
    total_ready_entries = '0;
    indv_rs_we = '0;
    for(int i = 0; i < RS_SIZE; i++) begin
        //this if condition is hella sus if it works thank god but idk
        if(indv_rs_write_rdy[i] == 1'b1 && rs_we[s] == 1'b1 && s < PIPE_WIDTH) begin
             rs_sel[i][s] = 1'b1;
             indv_rs_we[i] = 1'b1;
             s = s + 1'b1;
        end
        total_open_entries += indv_rs_write_rdy[i];
        total_ready_entries += indv_rs_read_rdy[i];
        muxed_rs_entry[i] = rs_entry[oh_2_i(rs_sel[i])];
    end
    for(int i = 0; i < PIPE_WIDTH; i++) rs_rdy[i] = (total_open_entries > i + 1) ? 1 : 0;

    //outputs
    c1 = ret_exe_candidate(1);
    c2 = ret_exe_candidate(2);
    foreach(execute_pkt[i]) execute_pkt[i] = '0;
    if(total_ready_entries > 0) begin
        if(^alu_rdy == 1'b1) begin
            indv_alu_rdy[c1] = 1'b1;
            if(alu_rdy[0]) execute_pkt[0] = indv_execute_pkt[c1];
            else execute_pkt[1] = indv_execute_pkt[c1];  
        end
        else if (alu_rdy == 2'b11 && total_ready_entries == 1) begin
            indv_alu_rdy[c1] = 1'b1;
            execute_pkt[0] = indv_execute_pkt[c1];

        end
        else if(alu_rdy == 2'b11) begin
            indv_alu_rdy[c1] = 1'b1;
            indv_alu_rdy[c2] = 1'b1;
            execute_pkt[0] = indv_execute_pkt[c1];
            execute_pkt[1] = indv_execute_pkt[c2];
        end
    end
end

//logic to select open reservation stations and write to them
//if possible  select lowest  2 reservation stations
//if 1 res station open and 2 entries, select entry 0, and flip flip_count, next time select entry 1 and flip...




endmodule