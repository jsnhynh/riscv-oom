`timescale 1ns/1ps
import riscv_isa_pkg::*;
import uarch_pkg::*;

module cpu_tb;

    //-------------------------------------------------------------
    // Test Configuration
    //-------------------------------------------------------------
    localparam TEST_FILE = "rv32im_test.hex";
    localparam MAX_CYCLES = 100000;

    //-------------------------------------------------------------
    // Test Statistics
    //-------------------------------------------------------------
    int tests_passed = 0;
    int tests_failed = 0;
    int assertions_checked = 0;
    int cycle_count = 0;
    int instruction_count = 0;
    real ipc;

    //-------------------------------------------------------------
    // Clock and Reset
    //-------------------------------------------------------------
    logic clk;
    logic rst;

    initial begin
        clk = 0;
        forever #(CLK_PERIOD/2) clk = ~clk;
    end

    //-------------------------------------------------------------
    // DUT Instantiation
    //-------------------------------------------------------------
    cpu #(
        .SIMPLE_MEM_MODE(1)
    ) dut (
        .clk(clk),
        .rst(rst)
    );

    //-------------------------------------------------------------
    // Instruction Tracking
    //-------------------------------------------------------------
    always_ff @(posedge clk) begin
        if (!rst) begin
            // Count committed instructions by monitoring ROB commit
            // Assumes commit_write_ports indicate valid commits
            for (int i = 0; i < PIPE_WIDTH; i++) begin
                if (dut.core0.commit_write_ports[i].we) begin
                    instruction_count++;
                end
            end
        end
    end

    //-------------------------------------------------------------
    // Helper Tasks
    //-------------------------------------------------------------
    
    task automatic check_assertion(
        input string test_name,
        input logic condition,
        input string fail_msg
    );
        assertions_checked++;
        if (condition) begin
            $display("  [PASS] %s", test_name);
            tests_passed++;
        end else begin
            $display("  [FAIL] %s: %s", test_name, fail_msg);
            tests_failed++;
        end
    endtask

    task automatic check_register(
        input string test_name,
        input int reg_num,
        input logic [31:0] expected_value
    );
        logic [31:0] actual_value;
        actual_value = dut.core0.rename_stage.prf.registers[reg_num];
        
        assertions_checked++;
        if (actual_value == expected_value) begin
            $display("  [PASS] %s: x%0d = 0x%08h", test_name, reg_num, actual_value);
            tests_passed++;
        end else begin
            $display("  [FAIL] %s: x%0d = 0x%08h (expected 0x%08h)", 
                     test_name, reg_num, actual_value, expected_value);
            tests_failed++;
        end
    endtask

    task automatic check_memory(
        input string test_name,
        input logic [31:0] addr,
        input logic [31:0] expected_value
    );
        logic [31:0] actual_value;
        logic [7:0] byte0, byte1, byte2, byte3;
        
        byte0 = dut.mem.dmem[addr + 0];
        byte1 = dut.mem.dmem[addr + 1];
        byte2 = dut.mem.dmem[addr + 2];
        byte3 = dut.mem.dmem[addr + 3];
        actual_value = {byte3, byte2, byte1, byte0};
        
        assertions_checked++;
        if (actual_value == expected_value) begin
            $display("  [PASS] %s: mem[0x%h] = 0x%08h", test_name, addr, actual_value);
            tests_passed++;
        end else begin
            $display("  [FAIL] %s: mem[0x%h] = 0x%08h (expected 0x%08h)",
                     test_name, addr, actual_value, expected_value);
            tests_failed++;
        end
    endtask

    task automatic wait_for_completion();
        logic [31:0] completion_reg;
        logic done;
        int last_inst_count;
        int stall_cycles;
        
        done = 0;
        cycle_count = 0;
        stall_cycles = 0;
        last_inst_count = 0;
        
        $display("\n[INFO] Waiting for program completion (x31 = 0xFF or timeout)...\n");
        
        while (!done && cycle_count < MAX_CYCLES) begin
            @(posedge clk);
            cycle_count++;
            
            completion_reg = dut.core0.rename_stage.prf.registers[31];
            
            if (completion_reg == 32'hFF) begin
                done = 1;
                $display("[INFO] Program completed after %0d cycles", cycle_count);
                $display("[INFO] Instructions committed: %0d", instruction_count);
                if (cycle_count > 0) begin
                    ipc = real'(instruction_count) / real'(cycle_count);
                    $display("[INFO] IPC: %0.3f\n", ipc);
                end
            end
            
            // Print progress every 100 cycles
            if (cycle_count % 100 == 0) begin
                int insts_this_period = instruction_count - last_inst_count;
                real period_ipc = real'(insts_this_period) / 100.0;
                $display("[INFO] Cycle %0d: Instructions=%0d (+%0d), IPC=%0.3f, x31=0x%08h", 
                         cycle_count, instruction_count, insts_this_period, period_ipc, completion_reg);
                last_inst_count = instruction_count;
            end
        end
        
        if (!done) begin
            $display("[WARNING] Program did not complete within %0d cycles", MAX_CYCLES);
            $display("[WARNING] Final instruction count: %0d\n", instruction_count);
        end
        
        // Wait a few more cycles for pipeline to settle
        repeat(10) @(posedge clk);
        cycle_count += 10;
    endtask

    task automatic dump_registers();
        $display("\n========================================");
        $display("  Register File State");
        $display("========================================");
        for (int i = 0; i < 32; i += 4) begin
            $display("  x%02d=0x%08h  x%02d=0x%08h  x%02d=0x%08h  x%02d=0x%08h",
                     i,   dut.core0.rename_stage.prf.registers[i],
                     i+1, dut.core0.rename_stage.prf.registers[i+1],
                     i+2, dut.core0.rename_stage.prf.registers[i+2],
                     i+3, dut.core0.rename_stage.prf.registers[i+3]);
        end
        $display("========================================\n");
    endtask

    task automatic dump_performance_stats();
        $display("\n========================================");
        $display("  Performance Statistics");
        $display("========================================");
        $display("  Total Cycles:           %0d", cycle_count);
        $display("  Instructions Committed: %0d", instruction_count);
        if (cycle_count > 0) begin
            ipc = real'(instruction_count) / real'(cycle_count);
            $display("  IPC (Instructions/Cycle): %0.3f", ipc);
            $display("  CPI (Cycles/Instruction): %0.3f", 1.0/ipc);
        end
        $display("========================================\n");
    endtask

    //-------------------------------------------------------------
    // Test Stimulus
    //-------------------------------------------------------------
    initial begin
        $dumpfile("cpu_tb.vcd");
        $dumpvars(0, cpu_tb);
        
        $display("========================================");
        $display("  RV32IM CPU Testbench Started");
        $display("========================================");
        $display("  Test Program: %s", TEST_FILE);
        $display("  Max Cycles: %0d", MAX_CYCLES);
        $display("========================================\n");
        
        // Reset
        rst = 1;
        repeat(5) @(posedge clk);
        rst = 0;
        
        // Wait for program to complete
        wait_for_completion();
        
        // Dump performance statistics
        dump_performance_stats();
        
        // Dump register file
        dump_registers();
        
        //-------------------------------------------------------------
        // Verify Results
        //-------------------------------------------------------------
        $display("[TEST VERIFICATION] Checking expected register values...\n");
        
        // Test 1: Basic Arithmetic
        $display("=== Test 1: Basic Arithmetic ===");
        check_register("ADD: 5 + 7", 3, 32'd12);
        check_register("SUB: 7 - 5", 4, 32'd2);
        
        // Test 2: Logical Operations
        $display("\n=== Test 2: Logical Operations ===");
        check_register("AND: 5 & 7", 5, 32'd5);
        check_register("OR: 5 | 7", 6, 32'd7);
        check_register("XOR: 5 ^ 7", 7, 32'd2);
        check_register("ANDI: 7 & 3", 8, 32'd3);
        check_register("ORI: 5 | 8", 9, 32'd13);
        check_register("XORI: 7 ^ 15", 10, 32'd8);
        
        // Test 3: Shifts
        $display("\n=== Test 3: Shift Operations ===");
        check_register("SLLI: 5 << 2", 11, 32'd20);
        check_register("SRLI: 7 >> 1", 12, 32'd3);
        check_register("SRAI: -8 >> 1", 14, 32'hFFFFFFFC);  // -4
        check_register("SLL: 5 << 7", 15, 32'd640);
        check_register("SRL: 7 >> 5", 16, 32'd0);
        check_register("SRA: -8 >> 5", 17, 32'hFFFFFFFF);  // -1
        
        // Test 4: Comparisons
        $display("\n=== Test 4: Comparison Operations ===");
        check_register("SLT: 5 < 7", 18, 32'd1);
        check_register("SLT: 7 < 5", 19, 32'd0);
        check_register("SLTU: 0xFFFFFFF8 < 5 (unsigned)", 20, 32'd0);
        check_register("SLTI: 5 < 10", 21, 32'd1);
        check_register("SLTIU: 5 < 3", 22, 32'd0);
        
        // Test 5: Upper Immediates
        $display("\n=== Test 5: Upper Immediate Operations ===");
        check_register("LUI: 0x12345000", 23, 32'h12345000);
        check_assertion("AUIPC executed", 
                       dut.core0.rename_stage.prf.registers[24] != 32'h0,
                       "AUIPC result is zero");
        
        // Test 6: Branches
        $display("\n=== Test 6: Branch Operations ===");
        check_register("Branches executed correctly", 25, 32'd5);
        
        // Test 7: JAL/JALR
        $display("\n=== Test 7: JAL/JALR Operations ===");
        check_register("JAL/JALR path completed", 25, 32'd5);
        check_assertion("JAL stored return address",
                       dut.core0.rename_stage.prf.registers[26] != 32'h0,
                       "Return address is zero");
        
        // Test 8: Multiply/Divide
        $display("\n=== Test 8: Multiply/Divide Operations (M extension) ===");
        check_register("MUL: 6 * 7", 3, 32'd42);
        check_register("MUL: 100 * 10", 6, 32'd1000);
        check_register("DIV: 100 / 10", 7, 32'd10);
        check_register("REM: 100 % 10", 8, 32'd0);
        check_register("MUL: 6 * -3 (negative)", 10, 32'hFFFFFFEE);  // -18
        
        // Test 9: Memory Operations
        $display("\n=== Test 9: Memory Operations ===");
        check_register("LW: Load word (42)", 11, 32'd42);
        check_register("LW: Load word (1000)", 12, 32'd1000);
        check_register("LW: Load word (10)", 13, 32'd10);
        check_register("LBU: Load unsigned byte", 15, 32'hAB);
        check_register("LB: Load signed byte", 16, 32'hFFFFFFAB);
        check_register("LHU: Load unsigned halfword", 18, 32'h1234);
        check_register("LH: Load signed halfword", 19, 32'h1234);
        check_memory("SW: Store word (42)", 32'h100, 32'd42);
        check_memory("SW: Store word (1000)", 32'h104, 32'd1000);
        check_memory("SW: Store word (10)", 32'h108, 32'd10);
        
        // Completion marker
        $display("\n=== Completion Check ===");
        check_register("Completion marker", 31, 32'hFF);
        
        //-------------------------------------------------------------
        // Final Performance Report
        //-------------------------------------------------------------
        dump_performance_stats();
        
        //-------------------------------------------------------------
        // Test Summary
        //-------------------------------------------------------------
        $display("\n========================================");
        $display("  Test Summary");
        $display("========================================");
        $display("  Execution Cycles:     %0d", cycle_count);
        $display("  Instructions Retired: %0d", instruction_count);
        if (cycle_count > 0) begin
            $display("  IPC:                  %0.3f", ipc);
        end
        $display("  Tests Passed:         %0d", tests_passed);
        $display("  Tests Failed:         %0d", tests_failed);
        $display("  Total Checks:         %0d", assertions_checked);
        $display("========================================");
        
        if (tests_failed == 0) begin
            $display("  ✓ ALL TESTS PASSED!");
        end else begin
            $display("  ✗ SOME TESTS FAILED!");
        end
        $display("========================================\n");
        
        if (tests_failed > 0) begin
            $fatal(1, "Test failures detected");
        end
        
        $finish;
    end

    //-------------------------------------------------------------
    // Timeout Watchdog
    //-------------------------------------------------------------
    initial begin
        #(MAX_CYCLES * CLK_PERIOD * 2);
        $display("\n[ERROR] Global testbench timeout!");
        $display("[ERROR] Cycles: %0d, Instructions: %0d", cycle_count, instruction_count);
        $finish;
    end

endmodule
