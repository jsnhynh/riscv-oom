import uarch_pkg::*;

